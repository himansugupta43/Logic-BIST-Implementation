module c432_1 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output reg N223,N329,N370,N421,N430,N431,N432;

reg N1_new, N4_new, N8_new, N11_new, N14_new, N17_new, N21_new, N24_new, N27_new, N30_new,
      N34_new, N37_new, N40_new, N43_new, N47_new, N50_new, N53_new, N56_new, N60_new, N63_new,
      N66_new, N69_new, N73_new, N76_new, N79_new, N82_new, N86_new, N89_new, N92_new, N95_new,
      N99_new, N102_new, N105_new, N108_new, N112_new, N115_new;


reg N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

initial begin
//Marker
end

always@(*) begin

N1_new = N1;
N4_new = N4;
N8_new = N8;
N11_new = N11;
N14_new = N14;
N17_new = N17;
N21_new = N21;
N24_new = N24;
N27_new = N27;
N30_new = N30;
N34_new = N34;
N37_new = N37;
N40_new = N40;
N43_new = N43;
N47_new = N47;
N50_new = N50;
N53_new = N53;
N56_new = N56;
N60_new = N60;
N63_new = N63;
N66_new = N66;
N69_new = N69;
N73_new = N73;
N76_new = N76;
N79_new = N79;
N82_new = N82;
N86_new = N86;
N89_new = N89;
N92_new = N92;
N95_new = N95;
N99_new = N99;
N102_new = N102;
N105_new = N105;
N108_new = N108;
N112_new = N112;
N115_new = N115;

N118=~N1_new;
N119=~N4_new;
N122=~N11_new;
N123=~N17_new;
N126=~N24_new;
N127=~N30_new;
N130=~N37_new;
N131=~N43_new;
N134=~N50_new;
N135=~N56_new;
N138=~N63_new;
N139=~N69_new;
N142=~N76_new;
N143=~N82_new;
N146=~N89_new;
N147=~N95_new;
N150=~N102_new;
N151=~N108_new;

N154=~(N118&N4_new);
N157=~(N8_new|N119);
N158=~(N14_new|N119);

N159=~(N122&N17_new);
N162=~(N126&N30_new);
N165=~(N130&N43_new);
N168=~(N134&N56_new);
N171=~(N138&N69_new);
N174=~(N142&N82_new);
N177=~(N146&N95_new);
N180=~(N150&N108_new);

N183=~(N21_new|N123);
N184=~(N27_new|N123);
N185=~(N34_new|N127);
N186=~(N40_new|N127);
N187=~(N47_new|N131);
N188=~(N53_new|N131);
N189=~(N60_new|N135);
N190=~(N66_new|N135);
N191=~(N73_new|N139);
N192=~(N79_new|N139);
N193=~(N86_new|N143);
N194=~(N92_new|N143);
N195=~(N99_new|N147);
N196=~(N105_new|N147);
N197=~(N112_new|N151);
N198=~(N115_new|N151);

N199=N154&N159&N162&N165&N168&N171&N174&N177&N180;

N203=~N199;
N213=~N199;
N223=~N199;

N224=N203^N154;
N227=N203^N159;
N230=N203^N162;
N233=N203^N165;
N236=N203^N168;
N239=N203^N171;

N242=~(N1_new&N213);
N243=N203^N174;
N246=~(N213&N11_new);
N247=N203^N177;
N250=~(N213&N24_new);
N251=N203^N180;

N254=~(N213&N37_new);
N255=~(N213&N50_new);
N256=~(N213&N63_new);
N257=~(N213&N76_new);
N258=~(N213&N89_new);
N259=~(N213&N102_new);
N260=~(N224&N157);
N263=~(N224&N158);
N264=~(N227&N183);
N267=~(N230&N185);
N270=~(N233&N187);
N273=~(N236&N189);
N276=~(N239&N191);
N279=~(N243&N193);
N282=~(N247&N195);
N285=~(N251&N197);
N288=~(N227&N184);
N289=~(N230&N186);
N290=~(N233&N188);
N291=~(N236&N190);
N292=~(N239&N192);
N293=~(N243&N194);
N294=~(N247&N196);
N295=~(N251&N198);

N296=N260&N264&N267&N270&N273&N276&N279&N282&N285;

N300=~N263;
N301=~N288;
N302=~N289;
N303=~N290;
N304=~N291;
N305=~N292;
N306=~N293;
N307=~N294;
N308=~N295;
N309=~N296;
N319=~N296;
N329=~N296;

N330=N309^N260;
N331=N309^N264;
N332=N309^N267;
N333=N309^N270;

N334=~(N8_new&N319);
N335=N309^N273;
N336=~(N319&N21_new);
N337=N309^N276;
N338=~(N319&N34_new);
N339=N309^N279;
N340=~(N319&N47_new);
N341=N309^N282;
N342=~(N319&N60_new);
N343=N309^N285;

N344=~(N319&N73_new);
N345=~(N319&N86_new);
N346=~(N319&N99_new);
N347=~(N319&N112_new);
N348=~(N330&N300);
N349=~(N331&N301);
N350=~(N332&N302);
N351=~(N333&N303);
N352=~(N335&N304);
N353=~(N337&N305);
N354=~(N339&N306);
N355=~(N341&N307);
N356=~(N343&N308);

N357=N348&N349&N350&N351&N352&N353&N354&N355&N356;

N360=~N357;
N370=~N357;

N371=~(N14_new&N360);
N372=~(N360&N27_new);
N373=~(N360&N40_new);
N374=~(N360&N53_new);
N375=~(N360&N66_new);
N376=~(N360&N79_new);
N377=~(N360&N92_new);
N378=~(N360&N105_new);
N379=~(N360&N115_new);

N380=~(N4_new&N242&N334&N371);
N381=~(N246&N336&N372&N17_new);
N386=~(N250&N338&N373&N30_new);
N393=~(N254&N340&N374&N43_new);
N399=~(N255&N342&N375&N56_new);
N404=~(N256&N344&N376&N69_new);
N407=~(N257&N345&N377&N82_new);
N411=~(N258&N346&N378&N95_new);
N414=~(N259&N347&N379&N108_new);

N415=~N380;

N416=N381&N386&N393&N399&N404&N407&N411&N414;

N417=~N393;
N418=~N404;
N419=~N407;
N420=~N411;

N421=~(N415|N416);

N422=~(N386&N417);

N425=~(N386&N393&N418&N399);

N428=~(N399&N393&N419);

N429=~(N386&N393&N407&N420);
N430=~(N381&N386&N422&N399);
N431=~(N381&N386&N425&N428);
N432=~(N381&N422&N425&N429);

end

endmodule