module bist_controller (
    input clk,    
    input [35:0] N,    
    input [3:0] s,    
    output reg [3:0] memory_s,
    output reg [35:0] memory_N,
    output reg found   
);

    reg [39:0] memory [0:63]; // (36-bit N + 4-bit value)
    integer i;
    reg [35:0] N_new;

    always@(negedge clk)
    begin
        N_new = N;
    end

    initial begin        

        found = 0;
        memory[0] = {36'b000000000000000000000000000000000000, 4'b0000};//0
        memory[1] = {36'b011110100111011110001010000101000000, 4'b1000};//8
        memory[2] = {36'b101011000111100100001110010111101101, 4'b1000};//7
        memory[3] = {36'b011011010101100000101010000101101000, 4'b0011};//4
        memory[4] = {36'b010110100011111001101010001101111000, 4'b0111};//9
        memory[5] = {36'b101001000100111000101001100010000000, 4'b1100};//9
        memory[6] = {36'b011111000001001100101111000000110010, 4'b1100};
        memory[7] = {36'b110100000011001000111100110000110000, 4'b0111};
        memory[8] = {36'b111010100110010100111110000000110000, 4'b1101};
        memory[9] = {36'b000001111100001100101010101111101000, 4'b0010};
        memory[10] = {36'b011110100001100000110010000000110000, 4'b1011};
        memory[11] = {36'b000000100000101001011111100100101000, 4'b0111};
        memory[12] = {36'b010011100101010110001000000111110000, 4'b0010};
        memory[13] = {36'b011111100111011100010010010101111101, 4'b0001};
        memory[14] = {36'b000010000000100100100110000111101000, 4'b1110};
        memory[15] = {36'b100111100100110111011101011110011000, 4'b0111};
        memory[16] = {36'b011010011011001001010101100101110000, 4'b1101};
        memory[17] = {36'b001101000000010100111001100001100010, 4'b0111};
        memory[18] = {36'b001010100101111100110010110111001000, 4'b1100};
        memory[19] = {36'b011010100110010100111000000000000110, 4'b0011};
        memory[20] = {36'b010100111110111000101111111111100000, 4'b0111};
        memory[21] = {36'b001111101001101000010111000111101000, 4'b1000};
        memory[22] = {36'b101010000001010001111101110011011000, 4'b0110};

    end

    always @(posedge clk) 
    begin
        found = 0;
        for (i = 0; i < 63; i = i + 1) 
        begin
            if (N_new == memory[i][39:4]) 
            begin
                memory_N = memory[i][39:4];
                memory_s = memory[i][3:0];
                if (s == memory[i][3:0]) 
                begin
                    found = 1;
                end 
            end
        end
    end
endmodule

